// need to write this later
